library IEEE;
use IEEE.std_logic_1164.all;

package I2c_pkg is
    type i2c_data_buf_t is array(0 to 7) of std_logic_vector(7 downto 0);
end I2c_pkg;


package body I2c_pkg is 
end package body I2c_pkg;